ReRAM Example

V1 TE 0 PWL (0 0 0.25u 1.8 0.5u 0 0.75u -1.8 1.0u 0.0)

XR0 TE 0 sky130_fd_pr_reram__reram_cell Tfilament_0=3.8e-9

.tran 0.1n 1.5u

.inc /foss/pdks/sky130B/libs.tech/ngspice/sky130_fd_pr_reram__reram_cell.spice

.control
set filetype=ascii
.endc

.end