ReRAM Example

.model sky130_fd_pr_reram__reram_model sky130_fd_pr_reram__reram_cell area_ox=0.1024e-12
+ area_ox = 0.1024e-12
+ Tox = 5.0
+ Tfilament_max = 4.9
+ Tfilament_min = 3.3
+ Eact_generation = 1.501
+ Eact_recombination  = 1.500
+ I_k1  = 6.140e-5
+ Tfilament_ref = 4.7249
+ V_ref = 0.430
+ velocity_k1 = 150
+ gamma_k0  = 16.5
+ gamma_k1  = -1.25 
+ Temperature_0 = 300
+ C_thermal = 3.1825e-16
+ tau_thermal = 0.23e-9
+ t_step  = 1.0e-9 
+ smoothing = 1e-7
+ Kclip = 200

V1 TE 0 PWL (0 0 0.25u 1.8 0.5u 0 0.75u -1.8 1.0u 0.0)

N1 TE 0 nFilament sky130_fd_pr_reram__reram_model

.tran 0.1n 1.5u

.ic v(nFilament)=3.8

.control
set filetype=ascii
pre_osdi /root/.volare/volare/sky130/versions/sky130B/libs.tech/ngspice/sky130_fd_pr_reram__reram_cell.osdi
run
.endc

.end
